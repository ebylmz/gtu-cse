`define CLOCK 4
`define DELAY 1250

module alu32_tb();

	reg [31:0] A, B;
	reg clk;
	reg [2:0]ALUop;
	wire [31:0] result;

	alu32 t(result, clk, A, B, ALUop);
	
	initial begin
		clk = 1'b0;

		// add
		ALUop = 3'b000; A = 32'b0000_0000_0000_0000_0000_0000_0000_1101; B = 32'b0000_0000_0000_0000_0000_0000_0000_1100;
		#`DELAY;

		ALUop = 3'b000; A = 32'b1000_0000_0000_0000_0000_0000_0000_1101; B = 32'b0000_0000_0000_0000_0000_0000_0101_1100;
		#`DELAY;
		
		// sub
		ALUop = 3'b001; A = 32'b0000_0000_0000_0000_0000_0000_0010_1101; B = 32'b0000_0000_0000_0000_0000_0000_0000_1111;
		#`DELAY;
		
		ALUop = 3'b001; A = 32'b1000_0000_0000_0000_0000_0000_0010_1101; B = 32'b0000_0000_0000_0000_0000_0000_0000_1111;
		#`DELAY;
		
		// mult
		ALUop = 3'b010; A = 32'b0000_0000_0000_0000_0000_0000_0000_0011; B = 32'b0000_0000_0000_0000_0000_0000_0000_0010;
		#`DELAY;
		
		// mult
		ALUop = 3'b010; A = 32'b0000_0000_0000_0000_0000_0000_0000_1111; B = 32'b0000_0000_0000_0000_0000_0000_0000_0101;
		#`DELAY;
		
		// xor
		ALUop = 3'b011; A = 32'b0000_0010_0000_0000_0000_0000_0000_1101; B = 32'b0000_0010_0000_0000_0000_0000_0000_1100;
		#`DELAY;
	
		// and
		ALUop = 3'b100; A = 32'b0000_0010_0000_0000_0000_0000_0000_1101; B = 32'b0000_0010_0000_0000_0000_0000_0000_1100;
		#`DELAY;
		
		// or
		ALUop = 3'b101; A = 32'b0000_0010_0000_0000_0000_0000_0000_1101; B = 32'b0000_0010_0000_0000_0000_0000_0000_1100;
		#`DELAY;
		
		//slt
		ALUop = 3'b110; A = 32'b0000_0010_0000_0000_0000_0000_0000_1111; B = 32'b0000_0010_0000_0000_0000_0000_0000_1100;
		#`DELAY;
	
		ALUop = 3'b110; A = 32'b0000_0010_0000_0000_0000_0000_0000_0101; B = 32'b0000_0010_0000_0000_0000_0000_0000_1100;
		#`DELAY;
		
		// nor
		ALUop = 3'b111; A = 32'b0000_0010_0000_0000_0000_0000_0000_1101; B = 32'b0000_0010_0000_0000_0000_0000_0000_1100;
		#`DELAY; $finish;

	end
	
	// define clock cycle
	always begin
		#4 clk = ~clk;
	end
		
	initial begin
		$monitor("time = %5d, ALUop = %3b, A = %32b, B = %32b, result = %32b", $time, ALUop, A, B, result);
	end
	
	

endmodule