module or32(Y, A, B);

	output[31:0] Y;
	input[31:0] A, B;
	
	or g31 (Y[31], A[31], B[31]);
	or g30 (Y[30], A[30], B[30]);
	or g29 (Y[29], A[29], B[29]);
	or g28 (Y[28], A[28], B[28]);
	
	or g27 (Y[27], A[27], B[27]);
	or g26 (Y[26], A[26], B[26]);
	or g25 (Y[25], A[25], B[25]);
	or g24 (Y[24], A[24], B[24]);
	
	or g23 (Y[23], A[23], B[23]);
	or g22 (Y[22], A[22], B[22]);
	or g21 (Y[21], A[21], B[21]);
	or g20 (Y[20], A[20], B[20]);
	
	or g19 (Y[19], A[19], B[19]);
	or g18 (Y[18], A[18], B[18]);
	or g17 (Y[17], A[17], B[17]);
	or g16 (Y[16], A[16], B[16]);
	
	or g15 (Y[15], A[15], B[15]);
	or g14 (Y[14], A[14], B[14]);
	or g13 (Y[13], A[13], B[13]);
	or g12 (Y[12], A[12], B[12]);
	
	or g11 (Y[11], A[11], B[11]);
	or g10 (Y[10], A[10], B[10]);
	or g9 (Y[9], A[9], B[9]);
	or g8 (Y[8], A[8], B[8]);
	
	or g7 (Y[7], A[7], B[7]);
	or g6 (Y[6], A[6], B[6]);
	or g5 (Y[5], A[5], B[5]);
	or g4 (Y[4], A[4], B[4]);
	
	or g3 (Y[3], A[3], B[3]);
	or g2 (Y[2], A[2], B[2]);
	or g1 (Y[1], A[1], B[1]);
	or g0 (Y[0], A[0], B[0]);

endmodule 